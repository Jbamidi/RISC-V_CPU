module imm_gen(input logic [31:0] instr, output logic [31:0] imm_out);

always_comb begin
    unique case(instr[6:0])
        //I-Type
        7'b0010011, 7'b0000011, 7'b1100111 : imm_out = {{20{instr[31]}},instr[31:20]};
        //S-Type
        7'b0100011: imm_out = {{20{instr[31]}},instr[31:25],instr[11:7]};
        //B-Type
        7'b1100011: imm_out = {{19{instr[31]}}, instr[31], instr[7], instr[30:25], instr[11:8], 1'b0};

        //U-Type
        7'b0110111, 7'b0010111: imm_out = {instr[31:12],12'b0};
        //J-type
        7'b1101111:imm_out = {{11{instr[31]}}, instr[31], instr[19:12], instr[20], instr[30:21], 1'b0};
        
        default: imm_out = 32'b0;



    endcase
end

endmodule